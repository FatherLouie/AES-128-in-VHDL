library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library work;
use work.Gates.all;
use work.muxes.all;

entity sbox is
	port (b: in std_logic_vector(7 downto 0); y: out std_logic_vector(7 downto 0));
end entity;

architecture struct of sbox is
type lookup is array (0 to 255) of std_logic_vector(7 downto 0);
signal l: lookup;
signal s: std_logic_vector(256*8 - 1 downto 0);
signal outp: std_logic_vector(7 downto 0);
begin
	l(0)<=x"63"; l(1)<=x"7c"; l(2)<=x"77"; l(3)<=x"7b"; l(4)<=x"f2"; l(5)<=x"6b"; l(6)<=x"6f"; l(7)<=x"c5";
	l(8)<=x"30"; l(9)<=x"01"; l(10)<=x"67"; l(11)<=x"2b"; l(12)<=x"fe"; l(13)<=x"d7"; l(14)<=x"ab"; l(15)<=x"76";
	l(16)<=x"ca"; l(17)<=x"82"; l(18)<=x"c9"; l(19)<=x"7d"; l(20)<=x"fa"; l(21)<=x"59"; l(22)<=x"47"; l(23)<=x"f0";
	l(24)<=x"ad"; l(25)<=x"d4"; l(26)<=x"a2"; l(27)<=x"af"; l(28)<=x"9c"; l(29)<=x"a4"; l(30)<=x"72"; l(31)<=x"c0";
	l(32)<=x"b7"; l(33)<=x"fd"; l(34)<=x"93"; l(35)<=x"26"; l(36)<=x"36"; l(37)<=x"3f"; l(38)<=x"f7"; l(39)<=x"cc";
	l(40)<=x"34"; l(41)<=x"a5"; l(42)<=x"e5"; l(43)<=x"f1"; l(44)<=x"71"; l(45)<=x"d8"; l(46)<=x"31"; l(47)<=x"15";
	l(48)<=x"04"; l(49)<=x"c7"; l(50)<=x"23"; l(51)<=x"c3"; l(52)<=x"18"; l(53)<=x"96"; l(54)<=x"05"; l(55)<=x"9a";
	l(56)<=x"12"; l(57)<=x"80"; l(58)<=x"d6"; l(59)<=x"e2"; l(60)<=x"eb"; l(61)<=x"27"; l(62)<=x"b2"; l(63)<=x"75";
	l(64)<=x"09"; l(65)<=x"83"; l(66)<=x"2c"; l(67)<=x"1a"; l(68)<=x"1b"; l(69)<=x"6e"; l(70)<=x"5a"; l(71)<=x"a0";
	l(72)<=x"52"; l(73)<=x"3b"; l(74)<=x"d6"; l(75)<=x"b3"; l(76)<=x"29"; l(77)<=x"e3"; l(78)<=x"2f"; l(79)<=x"84";
	l(80)<=x"53"; l(81)<=x"d1"; l(82)<=x"00"; l(83)<=x"ed"; l(84)<=x"20"; l(85)<=x"fc"; l(86)<=x"b1"; l(87)<=x"5b";
	l(88)<=x"6a"; l(89)<=x"cb"; l(90)<=x"be"; l(91)<=x"39"; l(92)<=x"4a"; l(93)<=x"4c"; l(94)<=x"58"; l(95)<=x"cf";
	l(96)<=x"d0"; l(97)<=x"ef"; l(98)<=x"aa"; l(99)<=x"fb"; l(100)<=x"43"; l(101)<=x"4d"; l(102)<=x"33"; l(103)<=x"85";
	l(104)<=x"45"; l(105)<=x"f9"; l(106)<=x"02"; l(107)<=x"7f"; l(108)<=x"50"; l(109)<=x"3c"; l(110)<=x"9f"; l(111)<=x"a8";
	l(112)<=x"51"; l(113)<=x"a3"; l(114)<=x"40"; l(115)<=x"8f"; l(116)<=x"92"; l(117)<=x"9d"; l(118)<=x"38"; l(119)<=x"f5";
	l(120)<=x"bc"; l(121)<=x"b6"; l(122)<=x"da"; l(123)<=x"21"; l(124)<=x"10"; l(125)<=x"ff"; l(126)<=x"f3"; l(127)<=x"d2";
	l(128)<=x"cd"; l(129)<=x"0c"; l(130)<=x"13"; l(131)<=x"ec"; l(132)<=x"5f"; l(133)<=x"97"; l(134)<=x"44"; l(135)<=x"17";
	l(136)<=x"c4"; l(137)<=x"a7"; l(138)<=x"7e"; l(139)<=x"3d"; l(140)<=x"64"; l(141)<=x"5d"; l(142)<=x"19"; l(143)<=x"73";
	l(144)<=x"60"; l(145)<=x"81"; l(146)<=x"4f"; l(147)<=x"dc"; l(148)<=x"22"; l(149)<=x"2a"; l(150)<=x"90"; l(151)<=x"88";
	l(152)<=x"46"; l(153)<=x"ee"; l(154)<=x"b8"; l(155)<=x"14"; l(156)<=x"de"; l(157)<=x"5e"; l(158)<=x"0b"; l(159)<=x"db";
	l(160)<=x"e0"; l(161)<=x"32"; l(162)<=x"3a"; l(163)<=x"0a"; l(164)<=x"49"; l(165)<=x"06"; l(166)<=x"24"; l(167)<=x"5c";
	l(168)<=x"c2"; l(169)<=x"d3"; l(170)<=x"ac"; l(171)<=x"62"; l(172)<=x"91"; l(173)<=x"95"; l(174)<=x"e4"; l(175)<=x"79";
	l(176)<=x"e7"; l(177)<=x"c8"; l(178)<=x"37"; l(179)<=x"6d"; l(180)<=x"8d"; l(181)<=x"d5"; l(182)<=x"4e"; l(183)<=x"a9";
	l(184)<=x"6c"; l(185)<=x"56"; l(186)<=x"f4"; l(187)<=x"ea"; l(188)<=x"65"; l(189)<=x"7a"; l(190)<=x"ae"; l(191)<=x"08";
	l(192)<=x"ba"; l(193)<=x"78"; l(194)<=x"25"; l(195)<=x"2e"; l(196)<=x"1c"; l(197)<=x"a6"; l(198)<=x"b4"; l(199)<=x"c6";
	l(200)<=x"e8"; l(201)<=x"dd"; l(202)<=x"74"; l(203)<=x"1f"; l(204)<=x"4b"; l(205)<=x"bd"; l(206)<=x"8b"; l(207)<=x"8a";
	l(208)<=x"70"; l(209)<=x"3e"; l(210)<=x"b5"; l(211)<=x"66"; l(212)<=x"48"; l(213)<=x"03"; l(214)<=x"f6"; l(215)<=x"0e";
	l(216)<=x"61"; l(217)<=x"35"; l(218)<=x"57"; l(219)<=x"b9"; l(220)<=x"86"; l(221)<=x"c1"; l(222)<=x"1d"; l(223)<=x"9e";
	l(224)<=x"e1"; l(225)<=x"f8"; l(226)<=x"98"; l(227)<=x"11"; l(228)<=x"69"; l(229)<=x"d9"; l(230)<=x"8e"; l(231)<=x"94";
	l(232)<=x"9b"; l(233)<=x"1e"; l(234)<=x"87"; l(235)<=x"e9"; l(236)<=x"ce"; l(237)<=x"55"; l(238)<=x"28"; l(239)<=x"df";
	l(240)<=x"8c"; l(241)<=x"a1"; l(242)<=x"89"; l(243)<=x"0d"; l(244)<=x"bf"; l(245)<=x"e6"; l(246)<=x"42"; l(247)<=x"68";
	l(248)<=x"41"; l(249)<=x"99"; l(250)<=x"2d"; l(251)<=x"0f"; l(252)<=x"b0"; l(253)<=x"54"; l(254)<=x"bb"; l(255)<=x"16";
	
--	reorg: process(l) is
--	begin
--		for i in 0 to 7 loop
--			for j in 0 to 255 loop
--				s(256*i + j) <= l(j)(i);
--			end loop;
--		end loop;
--	end process;	
--	
--	mux_logic: for k in 0 to 7 generate
--		mux: MUX_256x1 port map(i => s(256*k + 255 downto 256*k), s => b, y => outp(k));
--	end generate;
	
	outp <= l(to_integer(unsigned(b)));
	y <= outp;
end architecture;
